module extend(input [15:0] immediate,output [31:0] extened);
   assign extened = immediate;

endmodule // extend

     
