


module datamem(clk,MemWrite,MemRead,Addr,Wdata,Rdata);

	input clk;
	input [31:0] Addr;
	input MemWrite;
	input MemRead;
	input [31:0] Wdata;
	output reg [31:0] Rdata;

	reg [31:0] mem [31:0];	

	initial begin
		$readmemh("inputmem.hex", mem);
	end

	//memory write
	always@(posedge clk)
	begin
		if(MemWrite)
		begin
			$display("Writing %d -> Addr: %d",Wdata,Addr);
			mem[Addr] <= Wdata; 
		end

		if(MemRead)
			Rdata <= mem[Addr];
	end


endmodule
